ENTITY plausable IS
    PORT (
        GX : IN BIT;
        GXOK : OUT BIT
    );
END ENTITY;