entity twoscomplement is
    port (
        clk   : in std_logic;
        reset : in std_logic;
        
    );
end entity twoscomplement;

architecture behav of twoscomplement is

begin

    

end architecture;